*** SPICE deck for cell inverter{sch} from library inverter-assignment
*** Created on Wed Aug 16, 2023 17:38:30
*** Last revised on Wed Sep 06, 2023 17:48:37
*** Written on Wed Sep 06, 2023 17:48:50 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: inverter-assignment:inverter{sch}
Mnmos@0 OUT INP gnd gnd nmos L=0.022U W=0.176U
Mpmos@0 vdd INP OUT vdd pmos L=0.022U W=0.352U

* Spice Code nodes in cell cell 'inverter-assignment:inverter{sch}'
.include "G:\Acads\Sem 7\DIC\22nm_HP.pm"
v1 vdd gnd DC 0.8
v2 INP gnd pwl(0 0 100p 0.8 1n 0.8 1.1n 0 2n 0)
.tran 2.1n
.END
.END
